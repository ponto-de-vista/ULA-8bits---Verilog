module porta_not(A, S);
    input A;
    output S;

    assign S = ~A;
endmodule
